library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"37",X"37",X"7F",X"FF",X"EE",X"00",X"00",X"00",X"CE",X"CE",X"67",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"EE",X"FF",X"7F",X"37",X"37",X"7F",X"00",X"00",X"00",X"33",X"67",X"CE",X"CE",X"EF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"F0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"FF",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"EC",X"E8",X"C0",X"00",X"00",X"00",X"00",X"00",X"73",X"71",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E8",X"EC",X"00",X"00",X"00",X"00",X"00",X"30",X"71",X"73",
		X"EC",X"E8",X"C0",X"00",X"00",X"00",X"00",X"0F",X"73",X"71",X"30",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"0F",X"00",X"00",X"00",X"00",X"C0",X"E8",X"EC",X"0F",X"00",X"00",X"00",X"00",X"30",X"71",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"77",X"30",X"30",X"30",X"30",X"30",X"30",X"77",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"0F",X"0F",X"01",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"0F",X"0C",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",
		X"0F",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0C",
		X"0C",X"0C",X"0C",X"0F",X"0F",X"00",X"00",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",
		X"0F",X"00",X"00",X"0F",X"0F",X"0C",X"0C",X"0C",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"33",X"00",X"00",X"00",
		X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"07",X"0F",X"0F",
		X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"07",X"0F",X"0F",
		X"01",X"0B",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",
		X"01",X"01",X"0B",X"0F",X"0F",X"0B",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0B",X"01",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"01",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"00",
		X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0E",X"0C",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"0C",X"0E",X"07",X"03",X"03",X"07",X"0F",X"0F",
		X"06",X"06",X"0E",X"0E",X"0E",X"0E",X"06",X"06",X"0C",X"0C",X"0E",X"0F",X"0F",X"0E",X"0C",X"0C",
		X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"06",X"0F",X"0F",X"07",X"03",X"03",X"07",X"0E",X"0C",
		X"EE",X"FF",X"11",X"99",X"55",X"FF",X"EE",X"00",X"33",X"77",X"55",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",
		X"33",X"99",X"99",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"11",X"33",X"22",X"00",X"33",X"77",X"44",X"44",X"44",X"66",X"22",X"00",
		X"55",X"FF",X"FF",X"55",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"BB",X"AA",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"44",X"66",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"EE",X"FF",X"99",X"99",X"99",X"BB",X"22",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"11",X"22",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"44",X"00",
		X"88",X"88",X"88",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"77",X"33",X"11",X"00",X"00",
		X"99",X"AA",X"CC",X"FF",X"CC",X"AA",X"99",X"00",X"44",X"22",X"11",X"77",X"11",X"22",X"44",X"00",
		X"88",X"CC",X"EE",X"FF",X"88",X"88",X"88",X"00",X"00",X"11",X"33",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"44",X"22",X"11",X"00",X"44",X"22",X"11",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"15",X"15",X"19",X"22",X"CC",X"33",X"44",X"88",X"8A",X"8A",X"89",X"44",X"33",
		X"00",X"FF",X"FF",X"44",X"44",X"FF",X"FF",X"00",X"00",X"11",X"33",X"66",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"EE",X"FF",X"11",X"11",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"33",X"11",X"DD",X"99",X"FF",X"FF",X"11",X"00",X"66",X"44",X"55",X"44",X"77",X"77",X"44",X"00",
		X"00",X"00",X"CC",X"99",X"FF",X"FF",X"11",X"00",X"66",X"44",X"55",X"44",X"77",X"77",X"44",X"00",
		X"FF",X"FF",X"99",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"44",X"77",X"77",X"44",X"00",X"00",
		X"00",X"00",X"EE",X"FF",X"11",X"77",X"66",X"00",X"44",X"44",X"77",X"77",X"44",X"44",X"00",X"00",
		X"11",X"33",X"EE",X"CC",X"FF",X"FF",X"11",X"00",X"66",X"77",X"11",X"00",X"77",X"77",X"44",X"00",
		X"33",X"11",X"11",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"44",X"77",X"77",X"44",X"00",
		X"FF",X"FF",X"88",X"CC",X"88",X"FF",X"FF",X"00",X"77",X"77",X"33",X"11",X"33",X"77",X"77",X"00",
		X"FF",X"FF",X"CC",X"88",X"00",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"33",X"77",X"77",X"00",
		X"CC",X"EE",X"33",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"00",X"88",X"88",X"99",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"DD",X"EE",X"55",X"11",X"11",X"FF",X"EE",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"11",X"BB",X"EE",X"CC",X"FF",X"FF",X"11",X"00",X"33",X"77",X"44",X"44",X"77",X"77",X"44",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"BB",X"22",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",X"00",
		X"00",X"00",X"11",X"FF",X"FF",X"11",X"00",X"00",X"00",X"66",X"44",X"77",X"77",X"44",X"66",X"00",
		X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"88",X"CC",X"66",X"33",X"66",X"CC",X"88",X"00",X"77",X"77",X"00",X"00",X"00",X"77",X"77",X"00",
		X"CC",X"FF",X"33",X"EE",X"33",X"FF",X"CC",X"00",X"77",X"77",X"00",X"11",X"00",X"77",X"77",X"00",
		X"11",X"33",X"66",X"CC",X"66",X"33",X"11",X"00",X"44",X"66",X"33",X"11",X"33",X"66",X"44",X"00",
		X"00",X"00",X"99",X"FF",X"FF",X"99",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"77",X"77",X"00",
		X"33",X"11",X"99",X"99",X"DD",X"77",X"33",X"00",X"66",X"77",X"55",X"44",X"44",X"44",X"66",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0B",X"01",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"06",X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"08",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"06",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"0C",X"0C",X"0C",X"0E",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"00",X"03",X"02",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"19",X"00",X"0E",X"0B",X"09",X"0F",X"0E",X"00",X"07",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"00",X"77",X"33",X"3B",X"33",X"3B",X"37",X"37",X"0C",X"08",X"0C",X"07",X"0C",X"00",X"06",X"05",
		X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"66",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"04",X"06",X"02",X"03",X"00",X"0D",X"0C",X"0C",X"06",X"07",X"0F",X"0E",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0C",X"0E",X"07",X"0E",X"00",X"0E",X"0F",X"0F",
		X"FF",X"EE",X"CC",X"00",X"0E",X"0E",X"0C",X"00",X"CC",X"FF",X"33",X"00",X"01",X"0F",X"01",X"00",
		X"00",X"11",X"FF",X"66",X"22",X"AA",X"33",X"77",X"00",X"33",X"BB",X"BB",X"BB",X"33",X"00",X"88",
		X"EE",X"33",X"33",X"EE",X"00",X"11",X"33",X"EE",X"11",X"33",X"33",X"11",X"00",X"CC",X"FF",X"11",
		X"CC",X"EE",X"33",X"33",X"FF",X"11",X"00",X"CC",X"11",X"33",X"33",X"11",X"FF",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"FF",X"FF",
		X"FF",X"FF",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"F3",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F3",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"F0",
		X"F3",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"F0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"2F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"0F",X"8F",X"0F",X"1F",X"4F",X"0E",X"00",X"00",
		X"E1",X"61",X"43",X"43",X"81",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"43",X"43",X"C3",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"8E",X"0F",X"00",X"00",X"00",X"0C",X"0F",X"8F",X"0F",X"2F",
		X"FC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"F3",X"C0",X"00",X"00",X"00",X"00",
		X"D2",X"3B",X"3F",X"0C",X"08",X"00",X"00",X"00",X"30",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"6F",X"47",X"13",X"00",X"00",X"01",X"03",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"38",X"00",X"00",X"00",X"C0",X"C2",X"FF",X"FF",X"3C",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"30",X"30",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"17",X"7F",X"B7",X"43",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"CE",X"7F",X"EF",X"9E",X"78",X"F0",X"00",X"7F",X"FF",X"EF",X"FF",X"7F",X"87",X"F0",
		X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"77",X"00",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"F0",X"F4",X"60",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"60",X"78",X"F0",X"F4",X"60",X"00",
		X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"60",X"00",X"06",X"0D",X"0A",X"09",X"00",X"00",X"00",X"10",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"60",X"F0",X"00",X"00",X"00",X"30",X"70",X"7A",X"30",X"08",
		X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",
		X"40",X"22",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"20",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"8E",X"0E",X"27",X"03",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"2F",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0F",X"8F",X"2F",
		X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",
		X"B5",X"38",X"70",X"71",X"20",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"30",X"71",X"F7",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"00",X"00",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"00",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"EE",X"CC",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",
		X"F0",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"16",
		X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",
		X"E5",X"E5",X"E9",X"E9",X"E1",X"E9",X"01",X"00",X"F2",X"F2",X"F4",X"F4",X"F9",X"F4",X"00",X"00",
		X"00",X"F7",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"E9",X"E1",X"E9",X"E9",X"E5",X"00",X"00",X"00",X"F4",X"F9",X"F4",X"F4",X"F2",
		X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",X"00",
		X"77",X"FF",X"FF",X"FF",X"77",X"33",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"77",X"FF",X"FF",X"FF",X"F7",X"B7",X"00",X"00",X"00",X"20",X"30",X"30",X"10",X"07",
		X"00",X"00",X"00",X"88",X"EE",X"FF",X"FF",X"EE",X"00",X"88",X"EE",X"FF",X"F3",X"F3",X"FF",X"FF",
		X"2F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"0F",X"8F",X"0F",X"1F",X"4F",X"0E",X"00",X"00",
		X"E1",X"61",X"43",X"43",X"81",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"43",X"43",X"C3",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"8E",X"0F",X"00",X"00",X"00",X"0C",X"0F",X"8F",X"0F",X"2F",
		X"D2",X"3B",X"3F",X"0C",X"08",X"00",X"00",X"00",X"30",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",
		X"8E",X"0E",X"27",X"03",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"3C",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"0F",X"0F",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",
		X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FE",X"FC",X"F8",X"C0",X"00",X"00",
		X"E5",X"E5",X"E9",X"E9",X"E1",X"E9",X"01",X"00",X"F2",X"F2",X"F4",X"F4",X"F9",X"F4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"61",X"43",X"43",X"81",X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"3B",X"3F",X"0C",X"08",X"00",X"00",X"00",X"30",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"77",X"00",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"22",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"B5",X"38",X"70",X"71",X"20",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"F7",X"F7",X"F3",X"FF",X"FF",X"EC",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"11",X"00",
		X"00",X"F7",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"43",X"43",X"C3",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"10",
		X"00",X"00",X"00",X"00",X"0B",X"6F",X"47",X"13",X"00",X"00",X"01",X"03",X"03",X"01",X"01",X"01",
		X"00",X"01",X"17",X"7F",X"B7",X"43",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"10",
		X"00",X"30",X"60",X"00",X"06",X"0D",X"0A",X"09",X"00",X"00",X"00",X"10",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"20",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"2F",X"87",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"00",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",
		X"00",X"00",X"00",X"30",X"30",X"30",X"71",X"F7",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F7",X"00",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"8E",X"0F",X"00",X"00",X"00",X"0C",X"0F",X"8F",X"0F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"38",X"00",X"00",X"00",X"C0",X"C2",X"FF",X"FF",X"3C",
		X"00",X"0C",X"CE",X"7F",X"EF",X"9E",X"78",X"F0",X"00",X"7F",X"FF",X"EF",X"FF",X"7F",X"87",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"80",X"60",X"F0",X"00",X"00",X"00",X"30",X"70",X"7A",X"30",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0F",X"8F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",
		X"00",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"E8",X"00",X"00",X"00",X"00",X"77",X"FF",X"BF",X"3F",
		X"00",X"00",X"01",X"E9",X"E1",X"E9",X"E9",X"E5",X"00",X"00",X"00",X"F4",X"F9",X"F4",X"F4",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"EE",X"FF",X"FF",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"33",X"77",X"67",X"EF",X"FF",X"00",X"33",X"FF",X"FF",X"0F",X"09",X"09",X"0F",
		X"7F",X"7F",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"67",X"77",X"33",X"11",X"00",X"00",X"00",X"09",X"09",X"0F",X"FF",X"FF",X"33",X"00",X"00",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"77",X"77",X"FF",X"EF",X"EF",X"FF",X"33",X"FF",X"FF",X"FF",X"0F",X"09",X"09",X"0F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"FF",X"77",X"77",X"11",X"00",X"00",X"09",X"09",X"0F",X"FF",X"FF",X"FF",X"33",X"00",
		X"00",X"CC",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"77",X"FF",X"89",X"00",X"8F",X"00",X"00",X"77",X"FF",X"FF",X"1F",X"3F",X"7F",
		X"FF",X"FF",X"FF",X"EE",X"EE",X"CC",X"00",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"89",X"FF",X"FF",X"33",X"00",X"00",X"00",X"3F",X"1F",X"FF",X"FF",X"FF",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"67",X"67",X"67",X"77",X"77",
		X"FF",X"FF",X"1F",X"01",X"01",X"0F",X"9F",X"08",X"CC",X"CC",X"CC",X"CC",X"CC",X"EE",X"EE",X"6E",
		X"00",X"00",X"88",X"88",X"CC",X"EE",X"77",X"11",X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0F",X"8F",X"FF",X"33",X"00",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"FF",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"EF",X"EF",X"EF",X"FF",
		X"77",X"FF",X"FF",X"1F",X"01",X"01",X"0F",X"1F",X"CC",X"CC",X"88",X"88",X"CC",X"CC",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"EF",X"EF",X"77",X"77",X"33",X"11",X"00",
		X"01",X"01",X"0F",X"1F",X"FF",X"FF",X"FF",X"33",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"FF",X"FF",X"EF",X"EF",
		X"00",X"FF",X"8F",X"0C",X"0C",X"0F",X"09",X"09",X"FF",X"FF",X"7F",X"3F",X"3F",X"7F",X"7F",X"6E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"77",X"33",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"FF",X"FF",X"FF",X"33",X"11",X"00",X"EE",X"EE",X"CC",X"CC",X"CC",X"88",X"88",X"88",
		X"77",X"FF",X"FF",X"3F",X"19",X"19",X"19",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"67",X"EF",X"EF",X"FF",
		X"3F",X"19",X"19",X"19",X"3F",X"FF",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EF",X"67",X"67",X"33",X"11",X"00",X"00",
		X"CC",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",
		X"00",X"00",X"11",X"33",X"77",X"67",X"EF",X"FF",X"00",X"77",X"FF",X"FF",X"1F",X"01",X"01",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"FF",X"77",X"33",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"FF",X"77",X"33",X"00",X"00",X"00",X"01",X"01",X"1F",X"FF",X"FF",X"FF",X"11",X"00",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"11",X"33",X"33",X"77",X"77",X"77",X"77",
		X"77",X"FF",X"FF",X"CF",X"8E",X"8E",X"8E",X"CF",X"88",X"FF",X"FF",X"3F",X"17",X"17",X"17",X"3F",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"8E",X"8E",X"8E",X"CF",X"FF",X"FF",X"77",X"00",X"17",X"17",X"17",X"3F",X"FF",X"FF",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"FF",X"FF",X"FF",X"8F",X"0C",X"0C",X"8F",X"00",X"00",X"CC",X"FF",X"7F",X"3F",X"3F",X"7F",
		X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"77",X"77",X"77",X"FF",X"EE",X"00",
		X"0C",X"0C",X"8F",X"FF",X"FF",X"CC",X"00",X"00",X"3F",X"3F",X"7F",X"CC",X"00",X"00",X"00",X"00",
		X"A0",X"A0",X"A0",X"E2",X"70",X"62",X"62",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"70",X"62",X"60",X"20",X"20",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"70",X"F0",X"C0",X"F8",X"FC",X"00",X"00",X"00",X"00",X"30",X"70",X"D2",X"70",
		X"00",X"00",X"00",X"10",X"10",X"90",X"FC",X"FD",X"00",X"00",X"40",X"E0",X"00",X"F0",X"FF",X"FF",
		X"F8",X"C0",X"F0",X"70",X"10",X"00",X"00",X"00",X"D2",X"70",X"30",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"90",X"10",X"10",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"10",X"70",X"F0",X"C8",X"88",X"D0",X"70",X"30",X"30",X"30",X"34",X"F0",X"F0",X"70",
		X"00",X"00",X"10",X"30",X"73",X"F7",X"F7",X"F3",X"00",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"80",X"80",X"C0",X"40",X"40",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"D0",X"F0",X"F0",X"70",X"30",X"30",X"30",X"34",X"F0",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"77",X"F3",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",
		X"C0",X"80",X"C0",X"40",X"60",X"20",X"20",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"70",X"F0",X"C0",X"80",X"D0",X"70",X"30",X"30",X"30",X"34",X"F0",X"F0",X"70",
		X"00",X"00",X"10",X"30",X"70",X"F1",X"F0",X"F0",X"00",X"80",X"80",X"00",X"FF",X"FE",X"F0",X"F0",
		X"F0",X"B0",X"C0",X"60",X"20",X"30",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"80",X"80",X"00",X"00",X"00",X"00",
		X"11",X"60",X"00",X"00",X"02",X"00",X"91",X"C0",X"40",X"22",X"11",X"00",X"00",X"C0",X"30",X"88",
		X"42",X"13",X"21",X"10",X"55",X"55",X"77",X"00",X"20",X"00",X"CC",X"58",X"EC",X"44",X"54",X"00",
		X"60",X"00",X"C4",X"22",X"20",X"90",X"40",X"00",X"00",X"30",X"C0",X"10",X"22",X"66",X"44",X"00",
		X"00",X"D5",X"55",X"77",X"30",X"70",X"10",X"90",X"60",X"CC",X"44",X"C4",X"90",X"80",X"04",X"00",
		X"00",X"00",X"88",X"BB",X"99",X"99",X"F7",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"33",
		X"F7",X"99",X"99",X"BB",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"11",X"DD",X"AA",X"88",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"22",X"11",X"00",X"11",X"32",X"77",X"00",X"00",X"00",X"11",X"DD",X"FF",X"E6",X"CE",
		X"00",X"00",X"88",X"AA",X"DD",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",
		X"32",X"11",X"00",X"11",X"22",X"CC",X"00",X"00",X"E6",X"FF",X"DD",X"11",X"00",X"00",X"00",X"00",
		X"22",X"11",X"DD",X"AA",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"22",X"11",X"00",X"11",X"32",X"77",X"00",X"00",X"00",X"11",X"DD",X"FF",X"F7",X"DF",
		X"00",X"00",X"88",X"AA",X"DD",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",
		X"32",X"11",X"00",X"11",X"22",X"CC",X"00",X"00",X"F7",X"FF",X"DD",X"11",X"00",X"00",X"00",X"00",
		X"22",X"11",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",X"88",X"00",X"00",X"11",
		X"00",X"00",X"00",X"88",X"77",X"77",X"F9",X"FF",X"00",X"00",X"00",X"11",X"77",X"EE",X"CC",X"4C",
		X"00",X"00",X"00",X"88",X"EE",X"11",X"22",X"00",X"00",X"00",X"88",X"88",X"77",X"00",X"00",X"00",
		X"F9",X"77",X"77",X"88",X"00",X"00",X"00",X"00",X"CC",X"EE",X"77",X"11",X"00",X"00",X"00",X"00",
		X"00",X"44",X"AA",X"AA",X"DD",X"DD",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"66",X"22",X"11",X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"EE",X"FF",X"F3",X"EF",
		X"88",X"DD",X"DD",X"AA",X"AA",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"11",X"22",X"66",X"11",X"00",X"F3",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"DD",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"22",X"CC",X"44",X"00",
		X"00",X"00",X"00",X"CC",X"33",X"33",X"74",X"FF",X"00",X"00",X"00",X"11",X"BB",X"FF",X"EE",X"AE",
		X"00",X"00",X"00",X"AA",X"DD",X"11",X"11",X"00",X"44",X"CC",X"22",X"11",X"00",X"00",X"00",X"00",
		X"74",X"33",X"33",X"CC",X"00",X"00",X"00",X"00",X"EE",X"FF",X"BB",X"11",X"00",X"00",X"00",X"00",
		X"44",X"88",X"00",X"88",X"EE",X"11",X"00",X"88",X"EE",X"11",X"00",X"40",X"11",X"66",X"88",X"00",
		X"00",X"01",X"88",X"00",X"55",X"55",X"77",X"88",X"00",X"00",X"00",X"40",X"CC",X"44",X"CC",X"11",
		X"00",X"45",X"88",X"00",X"00",X"88",X"66",X"00",X"BB",X"66",X"00",X"00",X"22",X"44",X"88",X"00",
		X"00",X"55",X"55",X"77",X"00",X"22",X"11",X"11",X"22",X"CC",X"44",X"CC",X"00",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"27",X"27",X"12",
		X"07",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"27",X"27",X"02",X"00",X"00",X"00",
		X"00",X"07",X"07",X"03",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"7F",X"07",X"01",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"CF",X"2D",X"06",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"03",X"07",X"07",X"00",X"00",X"01",X"07",X"7F",X"0F",X"00",X"00",X"00",X"00",
		X"2D",X"CF",X"0C",X"08",X"00",X"00",X"00",X"00",X"0F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"03",X"0F",X"0F",X"0F",X"0F",X"03",X"27",X"37",X"17",X"03",X"01",X"00",X"00",
		X"00",X"08",X"08",X"08",X"8C",X"4F",X"2D",X"06",X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"03",X"07",X"07",X"00",X"00",X"00",X"01",X"03",X"17",X"37",X"27",X"03",X"00",
		X"2D",X"4F",X"8C",X"08",X"08",X"08",X"00",X"00",X"0F",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"C3",X"0F",X"0C",X"38",X"4B",X"0F",X"00",X"01",X"13",X"01",X"00",X"01",X"13",X"01",
		X"00",X"0F",X"DE",X"0F",X"12",X"0F",X"CE",X"0C",X"00",X"0C",X"1E",X"07",X"0F",X"0F",X"07",X"03",
		X"0F",X"0F",X"0F",X"06",X"0F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"0E",X"0E",X"0C",X"08",X"00",X"00",X"0D",X"00",X"30",X"61",X"C3",X"A7",X"4F",X"4E",X"6F",
		X"00",X"0F",X"4B",X"0D",X"4B",X"0F",X"03",X"01",X"10",X"30",X"69",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"1E",X"68",X"48",X"0C",X"0C",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"03",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"61",X"C3",X"87",X"0F",X"4E",X"6F",
		X"00",X"0C",X"86",X"0A",X"87",X"0F",X"03",X"01",X"00",X"06",X"86",X"86",X"0E",X"0C",X"0C",X"0C",
		X"30",X"F0",X"E0",X"08",X"0B",X"0F",X"07",X"00",X"3F",X"17",X"03",X"00",X"00",X"00",X"00",X"00",
		X"09",X"08",X"08",X"01",X"01",X"00",X"00",X"00",X"0E",X"1E",X"0F",X"0F",X"0F",X"0D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"61",X"C3",X"97",X"A7",X"2F",X"6F",
		X"0E",X"4B",X"0D",X"4B",X"0F",X"09",X"01",X"01",X"03",X"43",X"43",X"4B",X"0F",X"0E",X"0C",X"0C",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"07",X"0F",X"0F",X"06",X"2C",X"3C",X"1E",X"0F",X"0F",X"0F",X"03",X"03",
		X"00",X"00",X"10",X"F0",X"4B",X"0F",X"0C",X"00",X"00",X"70",X"E1",X"D3",X"37",X"6F",X"0F",X"00",
		X"C3",X"96",X"0F",X"9E",X"0B",X"08",X"01",X"01",X"08",X"0C",X"04",X"0E",X"0F",X"0F",X"0F",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",
		X"03",X"0B",X"0F",X"0F",X"0B",X"03",X"03",X"03",X"0E",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"02",X"05",X"00",X"00",X"00",X"03",X"0C",X"00",X"80",X"00",X"04",X"02",X"00",X"00",X"77",X"EE",
		X"08",X"19",X"04",X"00",X"07",X"04",X"04",X"00",X"80",X"01",X"03",X"00",X"0C",X"00",X"02",X"01",
		X"00",X"88",X"CC",X"22",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"04",X"08",
		X"00",X"07",X"04",X"04",X"00",X"00",X"11",X"11",X"00",X"0C",X"00",X"08",X"0C",X"02",X"89",X"01",
		X"00",X"00",X"00",X"06",X"08",X"03",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"4B",X"0F",X"01",X"03",X"08",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"0F",X"08",X"08",X"0A",X"0D",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"CC",X"0C",X"07",X"2D",X"03",X"07",X"0C",X"08",X"08",X"08",X"0F",X"0F",
		X"09",X"0A",X"08",X"0F",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",X"08",X"08",X"0C",X"07",X"03",X"00",
		X"00",X"00",X"01",X"07",X"0C",X"08",X"02",X"09",X"00",X"00",X"00",X"00",X"11",X"03",X"02",X"03",
		X"00",X"00",X"01",X"02",X"8B",X"09",X"0F",X"4B",X"00",X"08",X"0C",X"02",X"04",X"01",X"0F",X"0F",
		X"05",X"0A",X"0C",X"07",X"01",X"00",X"00",X"00",X"02",X"03",X"11",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"09",X"8B",X"02",X"01",X"00",X"00",X"00",X"0F",X"01",X"04",X"02",X"0C",X"08",X"00",X"00",
		X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"0D",X"00",X"01",X"01",X"25",X"07",X"07",X"23",X"33",
		X"00",X"0C",X"0C",X"1D",X"0F",X"0F",X"8B",X"89",X"33",X"23",X"67",X"CF",X"0E",X"01",X"0B",X"0E",
		X"07",X"08",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"08",X"08",X"04",X"03",X"00",X"0E",X"07",X"04",X"04",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"03",X"03",X"4B",X"0F",X"0F",
		X"0C",X"0E",X"02",X"0A",X"0A",X"0A",X"0F",X"0E",X"00",X"00",X"00",X"06",X"0E",X"08",X"08",X"07",
		X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"07",X"57",X"77",X"00",X"00",X"00",X"01",X"02",X"04",
		X"07",X"03",X"01",X"00",X"00",X"09",X"06",X"00",X"04",X"0C",X"0C",X"0E",X"0B",X"01",X"00",X"00",
		X"CC",X"8E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"03",X"03",X"11",X"11",X"00",
		X"0E",X"0E",X"0E",X"0F",X"0F",X"4D",X"CD",X"01",X"00",X"33",X"67",X"0F",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"88",X"00",X"00",X"00",X"08",X"08",X"04",X"03",X"00",
		X"01",X"03",X"03",X"02",X"04",X"08",X"00",X"00",X"0C",X"0C",X"0E",X"07",X"67",X"33",X"11",X"11",
		X"00",X"00",X"0F",X"03",X"00",X"0F",X"03",X"00",X"00",X"01",X"01",X"25",X"07",X"07",X"23",X"33",
		X"00",X"0C",X"0C",X"0C",X"0F",X"0F",X"8B",X"8B",X"00",X"00",X"07",X"0C",X"08",X"0F",X"08",X"08",
		X"08",X"0A",X"0E",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"08",
		X"07",X"07",X"07",X"03",X"03",X"09",X"06",X"00",X"0B",X"02",X"0E",X"0F",X"01",X"03",X"02",X"02",
		X"0C",X"0C",X"00",X"00",X"06",X"06",X"0C",X"02",X"00",X"03",X"03",X"4B",X"0F",X"0F",X"57",X"77",
		X"00",X"08",X"08",X"08",X"0F",X"0F",X"07",X"07",X"00",X"01",X"03",X"0E",X"0C",X"06",X"03",X"08",
		X"0E",X"00",X"00",X"08",X"0D",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"07",X"03",X"03",X"01",X"01",X"08",X"06",X"01",X"09",X"0B",X"0E",X"0F",X"00",X"0C",X"02",X"0C",
		X"00",X"00",X"06",X"03",X"06",X"0C",X"08",X"09",X"00",X"00",X"00",X"01",X"03",X"0E",X"0D",X"01",
		X"00",X"00",X"00",X"0E",X"03",X"CD",X"0C",X"07",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"0F",
		X"0D",X"0D",X"0A",X"0C",X"06",X"03",X"06",X"00",X"01",X"01",X"0D",X"0E",X"03",X"01",X"00",X"00",
		X"2D",X"07",X"0C",X"CD",X"03",X"0E",X"00",X"00",X"0F",X"0F",X"08",X"08",X"00",X"00",X"00",X"00",
		X"03",X"02",X"0E",X"08",X"00",X"00",X"C4",X"30",X"22",X"01",X"01",X"80",X"C0",X"23",X"00",X"00",
		X"02",X"22",X"22",X"00",X"70",X"50",X"70",X"00",X"CC",X"88",X"00",X"01",X"C0",X"40",X"C0",X"22",
		X"00",X"00",X"00",X"06",X"11",X"80",X"08",X"00",X"00",X"66",X"88",X"01",X"06",X"08",X"00",X"11",
		X"CC",X"70",X"50",X"70",X"44",X"89",X"89",X"89",X"00",X"F3",X"40",X"C0",X"44",X"44",X"22",X"88",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"92",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"10",X"83",X"71",X"F0",
		X"92",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"03",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E1",X"E1",X"C0",X"C0",X"00",X"00",X"00",X"70",X"61",X"03",X"27",X"07",
		X"20",X"70",X"30",X"30",X"38",X"3C",X"52",X"D2",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"E1",X"E1",X"80",X"00",X"00",X"00",X"00",X"27",X"03",X"61",X"70",X"00",X"00",X"00",X"00",
		X"52",X"3C",X"38",X"30",X"30",X"70",X"20",X"00",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"E1",X"E1",X"C0",X"C0",X"00",X"00",X"00",X"70",X"21",X"03",X"27",X"07",
		X"10",X"30",X"30",X"30",X"38",X"3C",X"52",X"D2",X"00",X"80",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"E1",X"E1",X"80",X"00",X"00",X"00",X"00",X"27",X"03",X"21",X"70",X"00",X"00",X"00",X"00",
		X"52",X"3C",X"38",X"30",X"30",X"30",X"10",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"80",X"00",X"00",
		X"00",X"06",X"86",X"84",X"F0",X"F0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"03",X"30",X"74",X"3C",X"1E",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"F0",X"F0",X"C0",X"0C",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"60",X"90",X"80",X"40",X"F0",X"F0",X"F0",X"F0",X"70",X"B0",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"F0",X"F0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"03",X"30",X"74",X"3C",X"1E",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"C0",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"30",X"C0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"00",X"00",
		X"00",X"20",X"E0",X"E0",X"C0",X"C3",X"C3",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"03",X"30",X"74",X"3C",X"1E",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"C3",X"C3",X"C0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"90",X"A0",X"40",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"00",X"00",
		X"00",X"06",X"60",X"E0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"00",X"70",X"70",X"30",X"78",X"78",
		X"20",X"70",X"30",X"30",X"B0",X"F0",X"F0",X"F0",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"E0",X"E0",X"E0",X"60",X"06",X"00",X"00",X"78",X"30",X"70",X"70",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"B0",X"30",X"30",X"70",X"20",X"00",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"00",
		X"40",X"00",X"10",X"70",X"00",X"80",X"00",X"00",X"20",X"10",X"80",X"40",X"20",X"00",X"C0",X"02",
		X"04",X"00",X"A0",X"20",X"00",X"70",X"50",X"70",X"20",X"20",X"40",X"40",X"08",X"D0",X"00",X"01",
		X"E0",X"30",X"00",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"30",X"C0",X"10",X"10",X"10",X"20",
		X"0C",X"70",X"50",X"70",X"08",X"20",X"10",X"00",X"00",X"C0",X"00",X"10",X"08",X"20",X"10",X"10",
		X"00",X"00",X"07",X"0F",X"0D",X"01",X"03",X"0F",X"00",X"00",X"0E",X"0F",X"03",X"00",X"0C",X"0F",
		X"01",X"03",X"01",X"0C",X"0F",X"03",X"00",X"0C",X"08",X"0C",X"08",X"03",X"0F",X"0C",X"00",X"03",
		X"0C",X"01",X"0F",X"01",X"0E",X"00",X"0F",X"00",X"0B",X"08",X"07",X"00",X"0F",X"08",X"07",X"00",
		X"0F",X"03",X"08",X"07",X"00",X"0F",X"00",X"0F",X"0F",X"0C",X"01",X"0E",X"00",X"0F",X"00",X"0F",
		X"0F",X"0F",X"00",X"07",X"0C",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"07",X"03",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"06",X"0C",X"07",X"03",X"07",X"00",X"01",X"03",
		X"00",X"00",X"00",X"0F",X"08",X"00",X"0E",X"03",X"00",X"11",X"00",X"0C",X"00",X"04",X"02",X"06",
		X"33",X"00",X"0C",X"0E",X"07",X"0F",X"0C",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"0C",X"00",X"0F",X"0C",X"08",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"77",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"01",X"0F",X"00",X"0F",X"0F",X"0F",
		X"08",X"0E",X"0F",X"0C",X"00",X"0E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"00",X"00",X"00",X"08",X"0C",X"0E",X"07",X"00",X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",X"0E",
		X"03",X"00",X"08",X"0C",X"0E",X"0F",X"0C",X"00",X"0E",X"0F",X"07",X"07",X"03",X"01",X"00",X"00",
		X"00",X"33",X"FF",X"EE",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"CC",
		X"00",X"77",X"77",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"11",X"00",X"88",X"00",X"33",
		X"FF",X"EE",X"88",X"00",X"0C",X"08",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"03",X"0F",X"03",X"00",X"FF",X"FF",X"FF",X"00",X"0F",X"0F",X"0E",X"00",
		X"88",X"CC",X"EE",X"EE",X"FF",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"33",X"77",X"77",X"33",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",
		X"CC",X"FF",X"FF",X"EE",X"88",X"33",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"33",
		X"33",X"77",X"77",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",
		X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",
		X"07",X"03",X"00",X"00",X"77",X"44",X"33",X"00",X"0F",X"0F",X"0F",X"00",X"22",X"99",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"BB",X"CC",X"44",X"66",X"33",X"22",X"33",
		X"77",X"44",X"FF",X"00",X"00",X"FF",X"77",X"00",X"EE",X"00",X"CC",X"00",X"00",X"EE",X"CC",X"00",
		X"03",X"01",X"00",X"08",X"0F",X"0F",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"01",X"00",
		X"07",X"0F",X"0C",X"08",X"08",X"0C",X"0E",X"0F",X"0E",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",
		X"0F",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0C",X"00",X"08",X"0C",X"0F",X"00",X"08",X"0F",X"0F",X"00",
		X"01",X"07",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"0E",X"08",X"00",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"0E",X"0F",X"0F",X"0E",X"0E",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0C",X"0F",X"0F",X"0C",X"0C",X"00",X"00",X"08",X"01",X"0F",X"0F",X"01",X"01",X"03",X"0F",
		X"00",X"00",X"08",X"0C",X"0C",X"0C",X"08",X"08",X"01",X"07",X"0E",X"0C",X"08",X"08",X"0C",X"0F",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0E",X"07",X"01",X"00",X"00",X"01",X"0F",
		X"0C",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"0F",X"00",X"00",X"07",X"0F",X"0C",X"00",X"00",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"0F",X"03",X"07");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
